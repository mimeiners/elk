* This models a jumper with series resistance of 1uOhm
.SUBCKT myjumper 1 2 3 4 5 6 7 8
.param j=limit(jres,1e-6,1e9)
R1 1 2 1e9
R2 3 4 1e9
R3 5 6 1e9
R4 7 8 1e-6
.ENDS
