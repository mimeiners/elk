* Motorola
* Semiconductor Databook (mid 1970s)
* 03 Jun 91	pwt	creation
.model D1N4001 D (Is=14.11n N=1.984 Rs=33.89m Ikf=94.81 Xti=3 Eg=1.11
+                 Cjo=25.89p M=.44 Vj=.3245 Fc=.5 Bv=75 Ibv=10u Tt=5.7u)
