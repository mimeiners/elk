*** Switching Diodes ***
.model D1N4148 D (Is=2.682n N=1.836 Rs=.5664 Ikf=44.17m Xti=3 Eg=1.11
+                 Cjo=4p M=.3333 Vj=.5 Fc=.5 Isr=1.565n Nr=2 Bv=100 Ibv=100u Tt=11.54n)
